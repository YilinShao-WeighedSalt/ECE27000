/home/shay/a/ece270/etc/lab11/tb_ll.sv